�P  ҄� �    @       @       @    @       @       @    @       @       @                             � � � �� � � �� �  �     0  �     0  �                                >  � � � >  � � � >  � ��� _����� _����� �   8  � �   8  � �                                �� � � �� � � �� ��7�������7�������7���  8p ���  8p ���          �        �     �� � � �� � � �� ��g�������g�������g��  pp��  pp��       p �     p �     ����� ?� ����� ?� ������O��?�����O��?�����O��<@�q��<@�q��<@        �        �     ����� ?� ����� ?� ����3�����?���3�����?���3����� <  � �� <  � �� <                               ����� ?� ����� ?� ����3�����?���3�����?���3������> `����> `����> `                             ���� � ���� � �����G������G������G��/�� "� ��/�� "� ��/��                               ���� � ���� � ���9��������9��������9�����'�8� �x��'�8� �x��'�8� �                             �� � � �� � � �� ��s�!���?���s�!���?���s� #�p�A�=�#�p�A�=�#�p�A�                             /� � � � /� � � � /� � �y�A�����y�A�����y�@��G���z���G���z���G��                               P @     P @     P \tAq��D\tAq��D\t@��#����?���#����?���#��                                                        � /@���� /@���� /@�/�0� ���/�0� ���/�0�                                                         ��� o������ o������     0  �     0  �                                                             ; � � N�; � � N�; �  �  @ 1  �  @ 1  �                                                             @       @       @    @       @       @    @       @       @                                @       @       @    @       @       @    @       @       @                                @       @       @    @       @       @    @       @       @                                @       @       @    @       @       @    @       @       @                                @       @       @    @       @       @    @       @       @                                @       @       @    @       @       @    @       @       @                                @       @       @    @       @       @    @       @       @                                @       @       @    @       @       @    @       @       @                                @       @       @    @       @       @    @       @       @                                @       @       @    @       @       @    @       @       @                                @       @       @    @       @       @    @       @       @                                @       @       @    @       @       @    @       @       @                                @       @       @    @       @       @    @       @       @                                @       @       @    @       @       @    @       @       @                                @       @       @    @       @       @    @       @       @                                @       @       @    @       @       @    @       @       @                                @       @       @    @       @       @    @       @       @                                                                                     ����������������������������                                                        �H �2Ֆ-�     �E� ��'����������������������������� ���?��*i����������3��+�                            �� ca�   @    �  �  `G�����������������������������8�����-����������A��'������                        �T7FA<&�P �    ��_�]��������������������������������ȹ���7�����������9=�٢@���                            �W�D�&Ȣ �  b�;-=��`�����������������������������Ǩ8�o��7]�������������� ��                           ��C6٤ �   ��ƃ��_���������������������������������n���&[��������g�39}��eW�                            ; \�� �&�i"1 `  
���;����������?����������?������ߣUr�m�q���������������P��                            ��"    � �      a � W���������������������������>W�������'�{��������������                            � *��	`9�@   C �f�,0 �W����������������������������� ���_���|�������������k�                                                                                     ���������������������������   @       @       @    @       @       @    @       @       @                                @       @       @    @       @       @    @       @       @                                @       @       @    @       @       @    @       @       @                                @       @       @    @       @       @    @       @       @                                @       @       @    @       @       @    @       @       @                                @       @       @    @       @       @    @       @       @                                @       @       @    @       @       @    @       @       @                                @       @       @    @       @       @    @       @       @                                @       @       @    @       @       @    @       @       @                                @       @       @    @       @       @    @       @       @                                @       @       @    @       @       @    @       @       @                                @       @       @    @       @       @    @       @       @                                @       @       @    @       @       @    @       @       @                                @       @       @    @       @       @    @       @       @                                @       @       @    @       @       @    @       @       @                                @       @       @    @       @       @    @       @       @                              �     0  �     0  �      @@   @@  � � � �� � � �� �                             �     ` �     ` �    @ @  @ @  @ ��� ������ ������        �        �     �  p a��  p a��   0��" � 0��" � 0���?��������?��������?��   p ��   p ��    p A�  p A�  `A�q�`A�q�`@��������������������  `p��  `p��    0p ��  0p ��   @   � @   � @ ��������������������0@�q�0@�q�0@    0  �     0  �     0  �     0  �     0  �  ?����������?����������?����� 0  � �  0  � �  0  �   8  � �   8  � �   0  �     0  �     0  �  ?����������?����������?����� 0 `��  0 `��  0 `�     ` �     ` �     @       @       @  ?����������?����������?�����. � "� ��. � "� ��. �  !� � �`!� � �`!� � �  ` �     ` �     `  ?����������?����������?�����  ``��  ``��  ` �@A  4 �@A  4 �@A  p !� �  p !� �  p  ?����������?����������?�����# 0� �0�# 0� �0�# 0� �k�A���k�A���k�A�  8 @�� 8 @�� 8 @���������������������  � `�  � `�  �   t � @   t � @   t  \ Ap� \ Ap� \ @����������������������#���.8���#���.8���#��     �        �        � @�= �� @�= �� @���?��������?��������?��/�� B��/�� B��/��        �        �     ��� O�?���� O�?���� ��� ������ ������       @       @                                 ; � � N�; � � N�; � � � � �� � � �� �  �  @ 1  �  @ 1  �     @       @       @    @       @       @    @       @       @                              �     0  �     0  �      @@   @@  � � � �� � � �� �                             �     ` �     ` �    @ @  @ @  @ ��� ������ ������        �        �     �  p a��  p a��   0��" � 0��" � 0���?��������?��������?��   p ��   p ��    p A�  p A�  `A�q�`A�q�`@��������������������  `p��  `p��    0p ��  0p ��   @   � @   � @ ��������������������0@�q�0@�q�0@    0  �     0  �     0  �     0  �     0  �  ?����������?����������?����� 0  � �  0  � �  0  �   8  � �   8  � �   0  �     0  �     0  �  ?����������?����������?����� 0 `��  0 `��  0 `�     ` �     ` �     @       @       @  ?����������?����������?�����. � "� ��. � "� ��. �  !� � �`!� � �`!� � �  ` �     ` �     `  ?����������?����������?�����  ``��  ``��  ` �@A  4 �@A  4 �@A  p !� �  p !� �  p  ?����������?����������?�����# 0� �0�# 0� �0�# 0� �k�A���k�A���k�A�  8 @�� 8 @�� 8 @���������������������  � `�  � `�  �   t � @   t � @   t  \ Ap� \ Ap� \ @����������������������#���.8���#���.8���#��     �        �        � @�= �� @�= �� @���?��������?��������?��/�� B��/�� B��/��        �        �     ��� O�?���� O�?���� ��� ������ ������       @       @                                 ; � � N�; � � N�; � � � � �� � � �� �  �  @ 1  �  @ 1  �     @       @       @    @       @       @    @       @       @                              �     0  �     0  �      @@   @@  � � � �� � � �� �                             �     ` �     ` �    @ @  @ @  @ ��� ������ ������        �        �     �  p a��  p a��   0��" � 0��" � 0���?��������?��������?��   p ��   p ��    p A�  p A�  `A�q�`A�q�`@��������������������  `p��  `p��    0p ��  0p ��   @   � @   � @ ��������������������0@�q�0@�q�0@    0  �     0  �     0  �     0  �     0  �  ?����������?����������?����� 0  � �  0  � �  0  �   8  � �   8  � �   0  �     0  �     0  �  ?����������?����������?����� 0 `��  0 `��  0 `�     ` �     ` �     @       @       @  ?����������?����������?�����. � "� ��. � "� ��. �  !� � �`!� � �`!� � �  ` �     ` �     `  ?����������?����������?�����  ``��  ``��  ` �@A  4 �@A  4 �@A  p !� �  p !� �  p  ?����������?����������?�����# 0� �0�# 0� �0�# 0� �k�A���k�A���k�A�  8 @�� 8 @�� 8 @���������������������  � `�  � `�  �   t � @   t � @   t  \ Ap� \ Ap� \ @����������������������#���.8���#���.8���#��     �        �        � @�= �� @�= �� @���?��������?��������?��/�� B��/�� B��/��        �        �     ��� O�?���� O�?���� ��� ������ ������       @       @                                 ; � � N�; � � N�; � � � � �� � � �� �  �  @ 1  �  @ 1  �     @       @       @    @       @       @    @       @       @                              �     0  �     0  �      @@   @@  � � � �� � � �� �                             �     ` �     ` �    @ @  @ @  @ ��� ������ ������        �        �     �  p a��  p a��   0��" � 0��" � 0���?��������?��������?��   p ��   p ��    p A�  p A�  `A�q�`A�q�`@��������������������  `p��  `p��    0p ��  0p ��   @   � @   � @ ��������������������0@�q�0@�q�0@    0  �     0  �     0  �     0  �     0  �  ?����������?����������?����� 0  � �  0  � �  0  �   8  � �   8  � �   0  �     0  �     0  �  ?����������?����������?����� 0 `��  0 `��  0 `�     ` �     ` �     @       @       @  ?����������?����������?�����. � "� ��. � "� ��. �  !� � �`!� � �`!� � �  ` �     ` �     `  ?����������?����������?�����  ``��  ``��  ` �@A  4 �@A  4 �@A  p !� �  p !� �  p  ?����������?����������?�����# 0� �0�# 0� �0�# 0� �k�A���k�A���k�A�  8 @�� 8 @�� 8 @���������������������  � `�  � `�  �   t � @   t � @   t  \ Ap� \ Ap� \ @����������������������#���.8���#���.8���#��     �        �        � @�= �� @�= �� @���?��������?��������?��/�� B��/�� B��/��        �        �     ��� O�?���� O�?���� ��� ������ ������       @       @                                 ; � � N�; � � N�; � � � � �� � � �� �  �  @ 1  �  @ 1  �     @       @       @    @       @       @    @       @       @                                                                                     ����������������������������                                                        ��;㎀ >�v���   V;����t�����������������������������?��q����?�������` |�                             ��� 5}��  /      .�@G������������������������������ �� �ʂ ?�����������J����                            �������  �B   ����?��������������������������������?`1���?���p�����U^?� `                               � p��=�c  � � /�����������������������������������������!'�������   �P                            �  8�� ]���   -j�����p��������������������������������eC���!�G����ҕ   �                            ���q%ZX��<�n�A@  ���w��?�`�����������������������������ڥ� ��p�����uw� ?� �                            O� � p�w�{���  F�Gw����`����������������������������?������ �H��n���x��    �                            �?��9����{����  W7c��  ����������������������������A�U�qr�DC?������Ȝ ?���                            �@ `^������ ,0T{�����0�����������������������������������
B"0�_����ϫ�D    �                            �> ���� ����   
 	@����P�������������������������������?�G	�B!���������   �                                                        @                           ����������������������������                                                                                                                                                                                                                                                             x � �   x � �   x �                              x � �   x � �   x �                              x � �   x � �   x �                              x � �   x � �   x �                              x � �   x � �   x �                              x � �   x � �   x �                              x � �   x � �   x �                              x � �   x � �   x �                              x � �   x � �   x �                              x � �   x � �   x �                              x � �   x � �   x �                              x � �   x � �   x �                              x � �   x � �   x �                              x � �   x � �   x �                              x � �   x � �   x �                              x � �   x � �   x �                              x � �   x � �   x �                              x � �   x � �   x �                              x � �   x � �   x �                              x � �   x � �   x �                              x � �   x � �   x �                              x � �   x � �   x �                              x � �   x � �   x �                              x � �   x � �   x �                              x � �   x � �   x �                              x � �   x � �   x �                              x � �   x � �   x �                              x � �   x � �   x �                              x � �   x � �   x �                              x � �   x � �   x �                              x � �   x � �   x �                              x � �   x � �   x �                              x � �   x � �   x �                              x � �   x � �   x �                              x � �   x � �   x �                              x � �   x � �   x �                             ����������������������������                            ����������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                 x � �   x � �   x �  x � �   x � �   x �  x � �   x � �   x �  x � �   x � �   x �  � 0 � 3  � 0 � 3  � 0  � 0 � 3  � 0 � 3  � 0  � 0 � 3  � 0 � 3  � 0  � 0 � 3  � 0 � 3  � 0  � 0 � 3  � 0 � 3  � 0  � 0 � 3  � 0 � 3  � 0  � 0 � 3  � 0 � 3  � 0  � 0 � 3  � 0 � 3  � 0  � 0 � 3  � 0 � 3  � 0  � 0 � 3  � 0 � 3  � 0  � 0 � 3  � 0 � 3  � 0  � 0 � 3  � 0 � 3  � 0  � 0 � 3  � 0 � 3  � 0  � 0 � 3  � 0 � 3  � 0  � 0 � 3  � 0 � 3  � 0  � 0 � 3  � 0 � 3  � 0  � 0 � 3  � 0 � 3  � 0  � 0 � 3  � 0 � 3  � 0  � 0 � 3  � 0 � 3  � 0  � 0 � 3  � 0 � 3  � 0  � 0 � 3  � 0 � 3  � 0  � 0 � 3  � 0 � 3  � 0  � 0 � 3  � 0 � 3  � 0  � 0 � 3  � 0 � 3  � 0  � 0 � 3  � 0 � 3  � 0  � 0 � 3  � 0 � 3  � 0  � 0 � 3  � 0 � 3  � 0  � 0 � 3  � 0 � 3  � 0  x � �   x � �   x �  x � �   x � �   x �  x � �   x � �   x �  x � �   x � �   x �                                                                                                                 d@         ���vy9�sN@�c�A���9`9�D�L�Y��	$�9��=gÎvsg,#�8�L'�<�7`���vy9�sN@�c�A���9`9�D�L�Y��	$�9��=gÎvsg,#�8�L'�<�7`                                                                  ���vy9�sN@�c�A���9`9�D�L�Y��	$�9��=gÎvsg,#�8�L'�<�7`�(QIEE"	�AAA�RA"��QE R�e$A	%YE%EH��QI�H� QR$AE����(QIEE"	�AAA�RA"��QE R�e$A	%YE%EH��QI�H� QR$AE���                                                                  �(QIEE"	�AAA�RA"��QE R�e$A	%YE%EH��QI�H� QR$AE����(IE}>	�OAAUA"��==�D�
H�E$BU�QE%�EO��I �H�C�=HDOE����(IE}>	�OAAUA"��==�D�
H�E$BU�QE%�EO��I �H�C�=HDOE���                                                                  �(IE}>	�OAAUA"��==�D�
H�E$BU�QE%�EO��I �H�C�=HDOE����(IEA 	�QAAUA"� EEPD@
D�E$BUQE%EH �I �H�DQEDDQE���(IEA 	�QAAUA"� EEPD@
D�E$BUQE%EH �I �H�DQEDDQE��                 P  @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @       �       �    0�?��  `@��  @ ��0@  �  ���0    �  ���0 `  @  ���  � �`  ��� `A p  ���� �A� 8 @�� � t \ @��#��   @�?���   � �      � �   @  @  @       �       �    0�?��  `@��  @ ��0@  �  ���0    �  ���0 `  @  ���  � �`  ��� `A p  ���� �A� 8 @�� � t \ @��#��   @�?���   � �      � �   @  @  @       �       �    0�?��  `@��  @ ��0@  �  ���0    �  ���0 `  @  ���  � �`  ��� `A p  ���� �A� 8 @�� � t \ @��#��   @�?���   � �      � �   @  @  @       �       �    0�?��  `@��  @ ��0@  �  ���0    �  ���0 `  @  ���  � �`  ��� `A p  ���� �A� 8 @�� � t \ @��#��   @�?���   � �      � �   @  @  @        x                                                                x                                                                                                                                  x                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 P    �       �    0�?��  `@��  @ ��0@  �  ���0    �  ���0 `  @  ���  � �`  ��� `A p  ���� �A� 8 @�� � t \ @��#��   @�?���   � �      � �   @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @       �       �    0�?��  `@��  @ ��0@  �  ���0    �  ���0 `  @  ���  � �`  ��� `A p  ���� �A� 8 @�� � t \ @��#��   @�?���   � �      � �   @  @  @       �       �    0�?��  `@��  @ ��0@  �  ���0    �  ���0 `  @  ���  � �`  ��� `A p  ���� �A� 8 @�� � t \ @��#��   @�?���   � �      � �   @  @  @       �       �    0�?��  `@��  @ ��0@  �  ���0    �  ���0 `  @  ���  � �`  ��� `A p  ���� �A� 8 @�� � t \ @��#��   @�?���   � �      � �   @  @  @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 P    �       �    0�?��  `@��  @ ��0@  �  ���0    �  ���0 `  @  ���  � �`  ��� `A p  ���� �A� 8 @�� � t \ @��#��   @�?���   � �      � �   @  @  @       �       �    0�?��  `@��  @ ��0@  �  ���0    �  ���0 `  @  ���  � �`  ��� `A p  ���� �A� 8 @�� � t \ @��#��   @�?���   � �      � �   @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @       �       �    0�?��  `@��  @ ��0@  �  ���0    �  ���0 `  @  ���  � �`  ��� `A p  ���� �A� 8 @�� � t \ @��#��   @�?���   � �      � �   @  @  @       �       �    0�?��  `@��  @ ��0@  �  ���0    �  ���0 `  @  ���  � �`  ��� `A p  ���� �A� 8 @�� � t \ @��#��   @�?���   � �      � �   @  @  @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 P    �       �    0�?��  `@��  @ ��0@  �  ���0    �  ���0 `  @  ���  � �`  ��� `A p  ���� �A� 8 @�� � t \ @��#��   @�?���   � �      � �   @  @  @       �       �    0�?��  `@��  @ ��0@  �  ���0    �  ���0 `  @  ���  � �`  ��� `A p  ���� �A� 8 @�� � t \ @��#��   @�?���   � �      � �   @  @  @       �       �    0�?��  `@��  @ ��0@  �  ���0    �  ���0 `  @  ���  � �`  ��� `A p  ���� �A� 8 @�� � t \ @��#��   @�?���   � �      � �   @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @       �       �    0�?��  `@��  @ ��0@  �  ���0    �  ���0 `  @  ���  � �`  ��� `A p  ���� �A� 8 @�� � t \ @��#��   @�?���   � �      � �   @  @  @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 P    �       �    0�?��  `@��  @ ��0@  �  ���0    �  ���0 `  @  ���  � �`  ��� `A p  ���� �A� 8 @�� � t \ @��#��   @�?���   � �      � �   @  @  @       �       �    0�?��  `@��  @ ��0@  �  ���0    �  ���0 `  @  ���  � �`  ��� `A p  ���� �A� 8 @�� � t \ @��#��   @�?���   � �      � �   @  @  @       �       �    0�?��  `@��  @ ��0@  �  ���0    �  ���0 `  @  ���  � �`  ��� `A p  ���� �A� 8 @�� � t \ @��#��   @�?���   � �      � �   @  @  @       �       �    0�?��  `@��  @ ��0@  �  ���0    �  ���0 `  @  ���  � �`  ��� `A p  ���� �A� 8 @�� � t \ @��#��   @�?���   � �      � �   @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 !  @  @  @    �       � �      � 7��   � g��   ��O��<@  �����<     �����> `   ��G���     ������ �   � s� �A�    � y�@G��    P \t@#��      /@�0�       �         �         @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     !  @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @     @  @  @    �       � �      � 7��   � g��   ��O��<@  �����<     �����> `   ��G���     ������ �   � s� �A�    � y�@G��    P \t@#��      /@�0�       �         �         @  @  @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      