�#                     ��|��|��|    �P�P�P    ���    ���    ������    � P� P� P    � P� P� P    �P�P�P    ������                                                      y
�y
�y
�   �
 �
 �
    �
 �
 �
    �
 �
 �
    �
 �
 �
    �
 �
 �
    �
 �
 �
    �
 �
 �
    x� x� x�                                                                                               ��|��|��|��|�P�P�P�P����������������� P� P� P� P� P� P� P� P�P�P�P�P��������                                                  y
�y
�y
�y
��
 �
 �
 �
 �
 �
 �
 �
 �
 �
 �
 �
 �
 �
 �
 �
 �
 �
 �
 �
 �
 �
 �
 �
 �
 �
 �
 �
 x� x� x� x�                                                                         