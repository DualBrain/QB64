�P   ˀ�                                                                                                         �                                                    �                                                                                                        �                                                    �                           �   x � �   x � �                                                    � �   x � �   x � �                          �                           �   x � �   x � �                                                    � �   x � �   x � �                          �                           � 3  � 0 � 3  � 0 � 3                                                   � � 3  � 0 � 3  � 0 � 3                         �                           � 3  � 0 � 3  � 0 � 3                                                   � � 3  � 0 � 3  � 0 � 3                         �                           � 3  � 0 � 3  � 0 � 3                                                   � � 3  � 0 � 3  � 0 � 3                         �                           � 3  � 0 � 3  � 0 � 3                                                   � � 3  � 0 � 3  � 0 � 3                         �                           � 3  � 0 � 3  � 0 � 3                                                   � � 3  � 0 � 3  � 0 � 3                         �                           � 3  � 0 � 3  � 0 � 3                                                   � � 3  � 0 � 3  � 0 � 3                         �                           � 3  � 0 � 3  � 0 � 3                                                   � � 3  � 0 � 3  � 0 � 3                         �                           � 3  � 0 � 3  � 0 � 3                                                   � � 3  � 0 � 3  � 0 � 3                         �                           � 3  � 0 � 3  � 0 � 3                                                   � � 3  � 0 � 3  � 0 � 3                         �                           � 3  � 0 � 3  � 0 � 3                                                   � � 3  � 0 � 3  � 0 � 3                         �                           � 3  � 0 � 3  � 0 � 3                                                   � � 3  � 0 � 3  � 0 � 3                         �                           � 3  � 0 � 3  � 0 � 3                                                   � � 3  � 0 � 3  � 0 � 3                         �                           � 3  � 0 � 3  � 0 � 3                                                   � � 3  � 0 � 3  � 0 � 3                         �                           � 3  � 0 � 3  � 0 � 3                                                   � � 3  � 0 � 3  � 0 � 3                         �                           �   x � �   x � �                                                    � �   x � �   x � �                          �                           �   x � �   x � �                                                    � �   x � �   x � �                          �                                                                                                        �                                                    �                                                                                                        �                                                    �                                                                                                        �                                                    �                                                                                                        �                                                    �                                                                                                        �                                                    �                                                                                                        �                                                    �                                                                                                        �                                                    �                                                                                                        �                                                    �                                                                                                        �������������������������������                       �                                                                                                        �������������������������������                       �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                      � �   �         � �   �        � �   �         � �   �         �                                                                                      � �   �         � �   �        � �   �         � �   �         �                                                                                     � �   �        � �   �        � �   �        � �   �         �                                                                                     � �   �        � �   �        � �   �        � �   �         �                                                                                     � �   � ��     � �   � ��     � �   ���     � �   � ��      �                                                                                     � �   � ��     � �   � ��     � �   ���     � �   � ��      �                                                                                     � �   � ��     � �   � ��     � �   ���     � �   � ��      �                                                                                     � �   � ��     � �   � ��     � �   ���     � �   � ��      �                                                                                     �����������     �����������     �����������     �����������      �                                                                                     �����������     �����������     �����������     �����������      �                                                                                     �����������     �����������     �����������     �����������      �                                                                                     �����������     �����������     �����������     �����������      �                                                                                     ����������<     ����������<     ����������x     ����������<      �                                                                                     ����������<     ����������<     ����������x     ����������<      �                                                                                     ����������<     ����������<     ?����������x     ����������<      �                                                                                     ����������<     ����������<     ?����������x     ����������<      �                                                                                     ?��?�� ���<    ?��?�� ���<    ��� ���x>    ?��?�� ���<     �                                                                                     ?��?�� ���<    ?��?�� ���<    ��� ���x>    ?��?�� ���<     �                                                                                     ?���� ���<?    ?���� ���<?    ǀ�� ���x~    ?���� ���<?     �                                                                                     ?���� ���<?    ?���� ���<?    ǀ�� ���x~    ?���� ���<?     �                                                                                     ���� ����<|    ���� ����<|    ����� ����x�    ���� ����<|     �                                                                                     ���� ����<|    ���� ����<|    ����� ����x�    ���� ����<|     �                                                                                     ����� ����<�    ����� ����<�   ���� ����y�    ����� ����<�     �                                                                                     ����� ����<�    ����� ����<�   ���� ����y�    ����� ����<�     �                                                                                     � �   ����?�    � �   ����?�   � �   �����    � �   ����?�     �                                                                                     � �   ����?�    � �   ����?�   � �   �����    � �   ����?�     �                                                                                     � �   ����?�    � �   ����?�   � �   �����    � �   ����?�     �                                                                                     � �   ����?�    � �   ����?�   � �   �����    � �   ����?�     �                                                                                     ������ ����    ������ ����   ������ ����    ������ ����     �                                                                                     ������ ����    ������ ����   ������ ����    ������ ����     �                                                                                     ������ ����    ������ ����   ������ ����    ������ ����     �                                                                                     ������ ����    ������ ����   ������ ����    ������ ����     �                                                                                      ����� ����        ����� ����       ���������        ����� ����        �                                                                                      ����� ����        ����� ����       ���������        ����� ����        �                                                                                      ����� ����        ����� ����       ���������        ����� ����        �                                                                                      ����� ����        ����� ����       ���������        ����� ����        �                                                                                      �   � �������     �   � �������    �  ��������     �   � �������     �                                                                                      �   � �������     �   � �������    �  ��������     �   � �������     �                                                                                      �   � �������     �   � �������    �  ��������     �   � �������     �                                                                                      �   � �������     �   � �������    �  ��������     �   � �������     �                                                                                      �   � ������     �   � ������    �  � ������     �   � ������     �                                                                                      �   � ������     �   � ������    �  � ������     �   � ������     �                                                                                      �   � ������     �   � ������    �  � ������     �   � ������     �                                                                                      �   � ������     �   � ������    �  � ������     �   � ������     �                                                                                      ����� ���<�     ����� ���<�    ����� ���x�     ����� ���<�     �                                                                                      ����� ���<�     ����� ���<�    ����� ���x�     ����� ���<�     �                                                                                      ����� ���<�     ����� ���<�    ����� ���x�     ����� ���<�     �                                                                                      ����� ���<�     ����� ���<�    ����� ���x�     ����� ���<�     �                                                                                      ����� ���?��     ����� ���?��    ����� �����     ����� ���?��     �                                                                                      ����� ���?��     ����� ���?��    ����� �����     ����� ���?��     �                                                                                      ����� ���?��     ����� ���?��    ����� ����      ����� ���?��     �                                                                                      ����� ���?��     ����� ���?��    ����� ����      ����� ���?��     �                                                                                      �   � ����      �   � ����     �  � ����      �   � ����      �                                                                                      �   � ����      �   � ����     �  � ����      �   � ����      �                                                                                      �   � ����      �   � ����     �  � ����      �   � ����      �                                                                                      �   � ����      �   � ����     �  � ����      �   � ����      �                                                                                      ����� ��?�      ����� ��?�     ����� ���      ����� ��?�      �                                                                                      ����� ��?�      ����� ��?�     ����� ���      ����� ��?�      �                                                                                      ����� ��?�      ����� ��?�     ����� ���      ����� ��?�      �                                                                                      ����� ��?�      ����� ��?�     ����� ���      ����� ��?�      �                                                                                      ����� �?����     ����� �?����    ����� ?�����     ����� �?����     �                                                                                      ����� �?����     ����� �?����    ����� ?�����     ����� �?����     �                                                                                      ����� ?�?����     ����� ?�?����    ����� �����     ����� ?�?����     �                                                                                      ����� ?�?����     ����� ?�?����    ����� �����     ����� ?�?����     �                                                                                      �   � ?�?���     �   � ?�?���    �  �  ���     �   � ?�?���     �                                                                                      �   � ?�?���     �   � ?�?���    �  �  ���     �   � ?�?���     �                                                                                      �   � ? ?���     �   � ? ?���    �  � ~ ���     �   � ? ?���     �                                                                                      �   � ? ?���     �   � ? ?���    �  � ~ ���     �   � ? ?���     �                                                                                      ����� ?           ����� ?          ����� ~           ����� ?           �                                                                                      ����� ?           ����� ?          ����� ~           ����� ?           �                                                                                      ����� >           ����� >          ����� |           ����� >           �                                                                                      ����� >           ����� >          ����� |           ����� >           �                                                                                      �����  �����      �����  �����     ����� �����      �����  �����      �                                                                                      �����  �����      �����  �����     ����� �����      �����  �����      �                                                                                      �����  �����      �����  �����     ����� �����      �����  �����      �                                                                                      �����  �����      �����  �����     ����� �����      �����  �����      �                                                                                       ��   �����       ��   �����      ��  �����       ��   �����      �                                                                                       ��   �����       ��   �����      ��  �����       ��   �����      �                                                                                       ��   �����       ��   �����      ��  �����       ��   �����      �                                                                                       ��   �����       ��   �����      ��  �����       ��   �����      �                                                                                       ��   � �       ��   � �      ��  ��       ��   � �      �                                                                                       ��   � �       ��   � �      ��  ��       ��   � �      �                                                                                       ��   � �       ��   � �      ��  ��       ��   � �      �                                                                                       ��   � �       ��   � �      ��  ��       ��   � �      �                                                                                    ������� � �    ������� � �    ���������    ������� � �      �                                                                                    ������� � �    ������� � �    ���������    ������� � �      �                                                                                    ������� � �    ������� � �    ���������    ������� � �      �                                                                                    ������� � �    ������� � �    ���������    ������� � �      �                                                                                    ������� � �    ������� � �    ���������    ������� � �      �                                                                                    ������� � �    ������� � �    ���������    ������� � �      �                                                                                    ������� � �    ������� � �    ���������    ������� � �      �                                                                                    ������� � �    ������� � �    ���������    ������� � �      �                                                                                      ��   � �      ��   � �      ��  ��      ��   � �      �                                                                                      ��   � �      ��   � �      ��  ��      ��   � �      �                                                                                      ��   � �      ��   � �      ��  ��      ��   � �      �                                                                                      ��   � �      ��   � �      ��  ��      ��   � �      �                                                                                      ��   � �      ��   � �      ��  ��      ��   � �      �                                                                                      ��   � �      ��   � �      ��  ��      ��   � �      �                                                                                      ��   � �      ��   � �      ��  ��      ��   � �      �                                                                                      ��   � �      ��   � �      ��  ��      ��   � �      �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �       >      @      @         @       !    A@                             >      @      @         @       !    A@                      �                                                                                      >      @      @         @       !    A@                      �              @@    @  @      @     H !         e �                            @@    @  @      @     H !         e �              �                                                                                             @@    @  @      @     H !         e �              �              @@    @  @      @     H !         � �                            @@    @  @      @     H !         � �              �                                                                                             @@    @  @      @     H !         � �              �        s�㝞NgE�Ӑ9`X�g&8Xx�0S,m�BI9�v8OY�0㝄����9	�8���              s�㝞NgE�Ӑ9`X�g&8Xx�0S,m�BI9�v8OY�0㝄����9	�8���      �                                                                                       s�㝞NgE�Ӑ9`X�g&8Xx�0S,m�BI9�v8OY�0㝄����9	�8���      �       <� ARQQH�E"�PE�e�H�)DdDQHT�IBIEQIDQR(�RD"�,�AE�QE#)$             <� ARQQH�E"�PE�e�H�)DdDQHT�IBIEQIDQR(�RD"�,�AE�QE#)$      �                                                                                      <� ARQQH�E"�PE�e�H�)DdDQHT�IBIEQIDQR(�RD"�,�AE�QE#)$      �        ��RQ_O�E"��EEPH�$|DD� �(I�U}QI|QS�!RH"�(��OA�|�)$              ��RQ_O�E"��EEPH�$|DD� �(I�U}QI|QS�!RH"�(��OA�|�)$      �                                                                                       ��RQ_O�E"��EEPH�$|DD� �(I�U}QI|QS�!RH"�(��OA�|�)$      �        �ARQPHE"�PEEPH�"@DE�(I�UAQI@QR!RH"�(�QAQ@B)$              �ARQPHE"�PEEPH�"@DE�(I�UAQI@QR!RH"�(�QAQ@B)$      �                                                                                       �ARQPHE"�PEEPH�"@DE�(I�UAQI@QR!RH"�(�QAQ@B)$      �        �ARQQH�M"�PEE H�iDDESH�I"EQIDQR(�RP"�(�QE4�QE")$              �ARQQH�M"�PEE H�iDDESH�I"EQIDQR(�RP"�(�QE4�QE")$      �                                                                                       �ARQQH�M"�PEE H�iDDESH�I"EQIDQR(�RP"�(�QE4�QE")$      �        r��^N'4���9D� '�8Dx�1$%�"9�NI9OQ��P �IȠ��8�!��8�%$              r��^N'4���9D� '�8Dx�1$%�"9�NI9OQ��P �IȠ��8�!��8�%$      �                                                                                       r��^N'4���9D� '�8Dx�1$%�"9�NI9OQ��P �IȠ��8�!��8�%$      �                                                                                                                                                    �                                                                                                                                                         �                                                                                                                                                          �                                                                                                                                                            �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                �������������������������������������������������������������������������������                                                                                �������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                              �������������������������������������������������������������������������������                                                                                �������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            