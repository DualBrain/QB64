�P   ˀ�                                                                                      �����������      ��                          �p    �����������      �                         ��                          ��                             �����������      ����������������������������?�    �����������      �                                 @       @                                   �����������      �@      @       @    �    �����������      �                         ��      @       @    ��                             �����������      ��                            p    �����������      �                           � �� � � �� � � �                               ����������<      �  0  �     0  �     0 �    ����������<      �                         ��                           ��                             ����������<      � � � >  � � � >  � � � 0    ����������<      �                           _����� _����� _��                               ����������<      |�8  � �   8  � �   8  � L�    ����������<      �                         ��                           ��                             ����������<       � � �� � � �� � �3p    ����������<      �                           �����7�������7�����                               ?��?�� ���<      8p ���  8p ���  8p ��      ?��?�� ���<     �                         ��    �        �        ���                             ?��?�� ���<     x�� � �� � � �� � ��    ?��?�� ���<     �                          �����g�������g�����                               ?���� ���<?     x�pp��  pp��  pp��E     ?���� ���<?     �                         �� p �     p �     p ���                             ?���� ���<?     P� ?� ����� ?� ����� ?�:�    ?���� ���<?     �                          ?�����O��?�����O��?���                               ���� ����<|       �q��<@�q��<@�q��      ���� ����<|     �                         ��    �        �        ���                             ���� ����<|     �� ?� ����� ?� ����� ?��    ���� ����<|     �                          ?���3�����?���3�����?���                               ����� ����<�     y�� �� <  � �� <  � ��      ����� ����<�     �                         ��                           ��                             ����� ����<�     P� ?� ����� ?� ����� ?��    ����� ����<�     �                          ?���3�����?���3�����?���                               � �   ����?�     �����> `����> `���     � �   ����?�     �                         ��                           ��                             � �   ����?�     yp� � ���� � ���� �|�    � �   ����?�     �                          ����G������G����                               � �   ����?�      � ��/�� "� ��/�� "� ��s@    � �   ����?�     �                         ��                           ��                             � �   ����?�     �� � ���� � ���� ��    � �   ����?�     �                          ���9��������9��������                               ������ ����     Rx��'�8� �x��'�8� �x��&@    ������ ����     �                         ��                           ��                             ������ ����     r�� � �� � � �� � �Y�    ������ ����     �                          ���?���s�!���?���s�!���?�                               ������ ����     v�=�#�p�A�=�#�p�A�=�L�    ������ ����     �                         ��                           ��                             ������ ����     	p� � /� � � � /� � � �30    ������ ����     �                          �����y�A�����y�A����                                ����� ����        Z��z���G���z���G���z��     ����� ����        �                         ��                           ��                              ����� ����        %P@     P @     P @  ~p     ����� ����        �                          q��D\tAq��D\tAq��D                                ����� ����          ��?���#����?���#����?��     ����� ����        �                         ��                           ��                              ����� ����        _�                           |P     ����� ����        �                           ��� /@���� /@���                                �   � �������     Z����/�0� ���/�0� ���      �   � �������     �                         ��                           ��                              �   � �������     %P                           y�     �   � �������     �                           o������ o������ o���                                �   � �������     v�0  �     0  �     0  �        �   � �������     �                         ��                           ��                              �   � �������     	P                           �     �   � �������     �                           � N�; � � N�; � � N�                                �   � ������     P@ 1  �  @ 1  �  @ 1 \@     �   � ������     �                         ��                           ��                              �   � ������     r�                           #�     �   � ������     �                                 @       @                                    �   � ������     {P      @       @           �   � ������     �                         ��      @       @    ��                              �   � ������     �                           _�     �   � ������     �                                 @       @                                    ����� ���<�     �      @       @     �     ����� ���<�     �                         ��      @       @    ��                              ����� ���<�     y0                                ����� ���<�     �                                 @       @                                    ����� ���<�     y�      @       @    m�     ����� ���<�     �                         ��      @       @    ��                              ����� ���<�     P                                ����� ���<�     �                                 @       @                                    ����� ���?��            @       @    [      ����� ���?��     �                         ��      @       @    ��                              ����� ���?��     �                           $�     ����� ���?��     �                                 @       @                                    ����� ���?��     x�      @       @           ����� ���?��     �                         ��      @       @    ��                              ����� ���?��     @                           �     ����� ���?��     �                                 @       @                                    �   � ����      p      @       @    L`     �   � ����      �                         ��      @       @    ��                              �   � ����      x�                           3�     �   � ����      �                                 @       @                                    �   � ����       p      @       @           �   � ����      �                         ��      @       @    ��                              �   � ����      �                           �     �   � ����      �                                 @       @                                    ����� ��?�      �      @       @           ����� ��?�      �                         ��      @       @    ��                              ����� ��?�      |p                           �     ����� ��?�      �                                 @       @                                    ����� ��?�       p      @       @    �     ����� ��?�      �                         ��      @       @    ��                              ����� ��?�      �                                 ����� ��?�      �                                 @       @                                    ����� �?����     �      @       @          ����� �?����     �                         ��      @       @    ��                              ����� �?����      p                           p�     ����� �?����     �                                 @       @                                    ����� ?�?����            @       @           ����� ?�?����     �                         ��      @       @    ��                              ����� ?�?����     �                           �     ����� ?�?����     �                                 @       @                                    �   � ?�?���     �      @       @     �     �   � ?�?���     �                         ��      @       @    ��                              �   � ?�?���      p                           0     �   � ?�?���     �                                 @       @                                    �   � ? ?���      �      @       @    c      �   � ? ?���     �                         ��      @       @    ��                              �   � ? ?���                                 �     �   � ? ?���     �                                 @       @                                    ����� ?                 @       @           ����� ?           �                         ��      @       @    ��                              ����� ?            �                           �     ����� ?           �                                 @       @                                    ����� >            �      @       @    b      ����� >           �                         ��      @       @    ��                              ����� >                                      �     ����� >           �                                 @       @                                    �����  �����      p      @       @          �����  �����      �                         ��      @       @    ��                              �����  �����      �                           b�     �����  �����      �                                @       @                                   �����  �����      ?�      @       @    �     �����  �����      �                         ��      @       @    ��                              �����  �����      F                                 �����  �����      �                                                                                      ��   �����      �                           ��      ��   �����      �                         �������������������������������                               ��   �����      �                           �      ��   �����      �                                                                                       ��   �����      ?� \ C-Yb�(     �d\� �B��      ��   �����      �                         �?�����������������������������                               ��   �����      �����Ҧ�/�������?ᛣ?����?�      ��   �����      �                          B                          H                                ��   � �      ?�� v0�m!       ;� � ���      ��   � �      �                         �������������������������������                               ��   � �      _s��������������������	��o�      ��   � �      �                                                                                   ��   � �      s��Ctd�l�     ��l%�e���{�`      ��   � �      �                         ������������������������������`                               ��   � �      ?�ʼ�����z���������?���$���      ��   � �      �                                                                                    ������� � �      ?��|tI�l�    �/���@� ��   ������� � �      �                         �������������������������������                            ������� � �      s�z������u����������M,=��	���p   ������� � �      �                          �                                                       ������� � �      ��~)1�m�@ �   !ɀ�h<������   ������� � �      �                         �������������������������������                            ������� � �      7��������e���������3���:U{�p   ������� � �      �                                                                                    ������� � �      3�ʨ�	"h� �    1�:� ng�   ������� � �      �                         �3�����?����������?����������g�                            ������� � �      ���5W-�ݗm���?�������_�����   ������� � �      �                          @                                                        ������� � �      ���"   ̀@      �@Eq��   ������� � �      �                         ����������������������������                            ������� � �      s������2������������`����o�   ������� � �      �                                                                                      ��   � �      ?�� B� ��4  0 2�h�  9E��     ��   � �      �                         �������������������������������                              ��   � �      O���U��i�g���������9��<��ƺ�?�     ��   � �      �                                                                                      ��   � �      6                            c`     ��   � �      �                         �0                           �`                              ��   � �      O�����������������������������     ��   � �      �                                 @       @                                    ��   � �      9�      @       @    |�     ��   � �      �                         ��      @       @    ��                              ��   � �      F                                 ��   � �      �                                 @       @                                    ��   � �      4       @       @           ��   � �      �                         ��      @       @    ��                              ��   � �      K�                           �     ��   � �      �                                 @       @                                                              @       @                             �                         ��      @       @    ��                                                �                           �                       �                                 @       @                                                      @       @       @    
�                       �                         ��      @       @    ��                                                ?�                           uP                       �                                 @       @                                                      :�      @       @    6�                       �                         ��      @       @    ��                                                E                            IP                       �                                 @       @                                                             @       @    `                       �                         ��      @       @    ��                                                ~�                           r�                       �                                 @       @                                                              @       @                             �                         ��      @       @    ��                                                �                           �                       �                                 @       @                                                      A�      @       @    �                       �                         ��      @       @    ��                                                >p                           zP                       �                                 @       @                                                              @       @    ;`                       �                         ��      @       @    ��                                                �                           D�                       �                                 @       @                                                              @       @    f�                       �                         ��      @       @    ��                                                �                           0                       �                                 @       @                                                      5       @       @    �                       �                         ��      @       @    ��                                                J�                           bP                       �                                 @       @                                                       �      @       @    `                        �                         ��      @       @    ��                                                p                           �                       �                                 @       @                                                      (      @       @                             �                         ��      @       @    ��                                                W�                           �                       �                                 @       @                                                              @       @    c                        �                         ��      @       @    ��                                                �                           �                       �                                 @       @                                                      @       @       @    �                       �                         ��      @       @    ��                                                ?�                           a                       �                                 @       @                                                       @      @       @    q�                       �                         ��      @       @    ��                                                �                                                  �                             0  �     0  �     0                                                     @@   @@   @@ `                       �                         ��� �� � � �� � � ���                                                }�                           �                       �                             ` �     ` �     `                                                     @  @ @  @ @  �                       �                         �������� ������ �����                                                �   �        �        �                        �                           p a��  p a��  p a�                                                  0 �" � 0��" � 0��" ��                       �                         ��������?��������?��������                                                O� p ��   p ��   p ��                        �                           p A�  p A�  p A�                                                   �q�`A�q�`A�q��                       �                         ������������������������                                                �`p��  `p��  `p��                        �                           0p ��  0p ��  0p ��                                                     � @   � @   �p                        �                         ������������������������                                                y��q�0@�q�0@�q��                       �                           0  �     0  �     0  �                                                    C    0  �     0  �     �                       �                         �������?����������?������������                                                �� �  0  � �  0  � � ~                       �                           8  � �   8  � �   8  �                                                   �    0  �     0  �     �                       �                         �������?����������?������������                                                }p��  0 `��  0 `��                         �                             ` �     ` �     `                                                   6      @       @     �                       �                         �������?����������?������������                                                I�� ��. � "� ��. � "� ��                        �                          `!� � �`!� � �`                                                  !�     ` �     ` �   �                       �                         �������?����������?������������                                                e�`��  ``��  ``��                        �                            4 �@A  4 �@A  4                                                   A� �  p !� �  p !� � �                       �                         �������?����������?������������                                                �0�# 0� �0�# 0� �0�                        �                          ��k�A���k�A���                                                   �� 8 @�� 8 @��x                        �                         ������������������������                                                f� `�  � `�  � `�                       �                           � @   t � @   t � @                                                  \!p� \ Ap� \ Ap�                         �                         ������������������������                                                #Ў.8���#���.8���#���.8��                       �                           �        �        �                                                     P= �� @�= �� @�= �                         �                         ��������?��������?��������                                                ~�B��/�� B��/�� B���                       �                              �        �        �                                                   ``O�?���� O�?���� O�?�?�                       �                         �������� ������ �����                                                �  @       @       @ @                       �                                                                                                         p� N�; � � N�; � � N�?�                       �                         ��� �� � � �� � � ���                                                �@ 1  �  @ 1  �  @ 1 @                       �                                 @       @                                                      ;       @       @                             �                         ��      @       @    ��                                                D�                           �                       �                             0  �     0  �     0                                                   [� @@   @@   @@~�                       �                         ��� �� � � �� � � ���                                                $p                                                  �                             ` �     ` �     `                                                     @  @ @  @ @ }@                       �                         �������� ������ �����                                                �   �        �        � �                       �                           p a��  p a��  p a�                                                  ` �" � 0��" � 0��" �~�                       �                         ��������?��������?��������                                                � p ��   p ��   p ��                       �                           p A�  p A�  p A�                                                  p�q�`A�q�`A�q�?�                       �                         ������������������������                                                �`p��  `p��  `p��@                       �                           0p ��  0p ��  0p ��                                                  3Q   � @   � @   ��                       �                         ������������������������                                                L��q�0@�q�0@�q�|p                       �                           0  �     0  �     0  �                                                   #    0  �     0  �                              �                         �������?����������?������������                                                r�� �  0  � �  0  � � �                       �                           8  � �   8  � �   8  �                                                   3    0  �     0  �     �                       �                         �������?����������?������������                                                q���  0 `��  0 `�� tp                       �                             ` �     ` �     `                                                   `�      @       @     �                       �                         �������?����������?������������                                                B� ��. � "� ��. � "� ��~0                       �                          `!� � �`!� � �`                                                  9��     ` �     ` �                           �                         �������?����������?������������                                                Fp`��  ``��  ``��g�                       �                            4 �@A  4 �@A  4                                                  @�� �  p !� �  p !� � m                        �                         �������?����������?������������                                                ?r0�# 0� �0�# 0� �0��                       �                          ��k�A���k�A���                                                   �� 8 @�� 8 @��@                       �                         ������������������������                                                q� `�  � `�  � `~�                       �                           � @   t � @   t � @                                                  `p� \ Ap� \ Ap�T�                       �                         ������������������������                                                ��.8���#���.8���#���.8�+P                       �                           �        �        �                                                     x�= �� @�= �� @�= �j                        �                         ��������?��������?��������                                                @B��/�� B��/�� B���                       �                              �        �        �                                                   p0O�?���� O�?���� O�?��                       �                         �������� ������ �����                                                �  @       @       @ }P                       �                                                                                                        �� N�; � � N�; � � N�                         �                         ��� �� � � �� � � ���                                                pp@ 1  �  @ 1  �  @ 1 _�                       �                                 @       @                                                      @       @       @    *�                       �                         ��      @       @    ��                                                ?�                           UP                       �                             0  �     0  �     0                                                   P @@   @@   @@
                        �                         ��� �� � � �� � � ���                                                 �                           u�                       �                             ` �     ` �     `                                                   x�@  @ @  @ @ U                        �                         �������� ������ �����                                                    �        �        � *�                       �                           p a��  p a��  p a�                                                  ��" � 0��" � 0��" �1                        �                         ��������?��������?��������                                                x0 p ��   p ��   p ��N�                       �                           p A�  p A�  p A�                                                   �q�`A�q�`A�q�M                        �                         ������������������������                                                �`p��  `p��  `p��2�                       �                           0p ��  0p ��  0p ��                                                  `   � @   � @   �                        �                         ������������������������                                                ��q�0@�q�0@�q�w�                       �                           0  �     0  �     0  �                                                   �    0  �     0  �                              �                         �������?����������?������������                                                 � �  0  � �  0  � � �                       �                           8  � �   8  � �   8  �                                                   �    0  �     0  �     �                       �                         �������?����������?������������                                                 0��  0 `��  0 `�� tP                       �                             ` �     ` �     `                                                          @       @      @                       �                         �������?����������?������������                                                �� ��. � "� ��. � "� ���                       �                          `!� � �`!� � �`                                                  ��     ` �     ` �                           �                         �������?����������?������������                                                 p`��  ``��  ``��q�                       �                            4 �@A  4 �@A  4                                                  �� �  p !� �  p !� � 0�                       �                         �������?����������?������������                                                 0�# 0� �0�# 0� �0�O                       �                          ��k�A���k�A���                                                  ��� 8 @�� 8 @��i�                       �                         ������������������������                                                 0 `�  � `�  � `0                       �                           � @   t � @   t � @                                                   1p� \ Ap� \ Ap��                       �                         ������������������������                                                ��.8���#���.8���#���.8�xp                       �                           �        �        �                                                       = �� @�= �� @�= �~                        �                         ��������?��������?��������                                                �B��/�� B��/�� B���                       �                              �        �        �                                                   �O�?���� O�?���� O�?�|�                       �                         �������� ������ �����                                                    @       @       @                        �                                                                                      � �   �         ~ � N�; � � N�; � � N��     � �   �         �                         ��� �� � � �� � � ���                              � �   �         �@ 1  �  @ 1  �  @ 1 |0     � �   �         �                                 @       @                                   � �   �         �      @       @    �    � �   �         �                         ��      @       @    ��                             � �   �                                      pP    � �   �         �                             0  �     0  �     0                                � �   � ��      � @@   @@   @@\     � �   � ��      �                         ��� �� � � �� � � ���                             � �   � ��                                   #�    � �   � ��      �                             ` �     ` �     `                                � �   � ��      @�@  @ @  @ @       � �   � ��      �                         �������� ������ �����                             � �   � ��      ?    �        �        � �    � �   � ��      �                           p a��  p a��  p a�                               �����������      ��" � 0��" � 0��" �}�    �����������      �                         ��������?��������?��������                             �����������         p ��   p ��   p ��p    �����������      �                           p A�  p A�  p A�                               �����������      �q�`A�q�`A�q�x`    �����������      �                         ������������������������                             �����������        `p��  `p��  `p���    �����������      �                           0p ��  0p ��  0p ��                               ����������<      �   � @   � @   ��    ����������<      �                         ������������������������                             ����������<        �q�0@�q�0@�q�|p    ����������<      �                           0  �     0  �     0  �                                ����������<      �    0  �     0  �     o`    ����������<      �                         �������?����������?������������                             ����������<        � �  0  � �  0  � � �    ����������<      �                           8  � �   8  � �   8  �                                ?��?�� ���<     �    0  �     0  �           ?��?�� ���<     �                         �������?����������?������������                             ?��?�� ���<       ��  0 `��  0 `�� �    ?��?�� ���<     �                             ` �     ` �     `                                ?���� ���<?     �      @       @     ]�    ?���� ���<?     �                         �������?����������?������������                             ?���� ���<?      � ��. � "� ��. � "� ��"P    ?���� ���<?     �                          `!� � �`!� � �`                               ���� ����<|     `�     ` �     ` �   ]     ���� ����<|     �                         �������?����������?������������                             ���� ����<|      `��  ``��  ``��"�    ���� ����<|     �                            4 �@A  4 �@A  4                               ����� ����<�     �� �  p !� �  p !� � <@    ����� ����<�     �                         �������?����������?������������                             ����� ����<�      0�# 0� �0�# 0� �0�C�    ����� ����<�     �                          ��k�A���k�A���                               � �   ����?�     ��� 8 @�� 8 @��1�    � �   ����?�     �                         ������������������������                             � �   ����?�        `�  � `�  � `NP    � �   ����?�     �                           � @   t � @   t � @                               � �   ����?�     �p� \ Ap� \ Ap�+�    � �   ����?�     �                         ������������������������                             � �   ����?�       �.8���#���.8���#���.8�TP    � �   ����?�     �                           �        �        �                                  ������ ����     �= �� @�= �� @�= ��    ������ ����     �                         ��������?��������?��������                             ������ ����       B��/�� B��/�� B��lP    ������ ����     �                              �        �        �                                ������ ����     �O�?���� O�?���� O�?�3�    ������ ����     �                         �������� ������ �����                             ������ ����         @       @       @ Lp    ������ ����     �                                                                                      ����� ����        ��� N�; � � N�; � � N�p�     ����� ����        �                         ��� �� � � �� � � ���                              ����� ����        � @ 1  �  @ 1  �  @ 1      ����� ����        �                                 @       @                                    ����� ����        �      @       @    �     ����� ����        �                         ��      @       @    ��                              ����� ����        ��                            0     ����� ����        �                                                       @                              �   � �������     ��                           ��     �   � �������     �                         �������������������������������                              �   � �������     �                            ~p     �   � �������     �                                                                                      �   � �������     � ?��8�  c�n�   `s����7M��     �   � �������     �                         �������������������������������                              �   � �������     ����\A����H���������F @Ȳ p     �   � �������     �                          �                                                           �   � ������     ����p�W��  �  �   �T~ ��     �   � ������     �                         �������������������������������                              �   � ������     �� ���� ���������������3p     �   � ������     �                                                                                      �   � ������     ��	��1� � � ��!   
�������     �   � ������     �                         �������������������������������                              �   � ������     ��������������U��|  f<p     �   � ������     �                                                                                      ����� ���<�     ��  H  `����F2   ����jS�     ����� ���<�     �                         �������������������������������                              ����� ���<�     ����������B| ���������   ��p     ����� ���<�     �                                                                                      ����� ���<�     ��@` ����� ����    ֯������     ����� ���<�     �                         �������������������������������                              ����� ���<�     ������qFQ?��"w�����)P�   �     ����� ���<�     �                                                                                      ����� ���?��     �O�U��=��v�x�   H��w����p     ����� ���?��     �                         �����������������������������p                              ����� ���?��     ����8�Zp�0�������Wp��� 	_�     ����� ���?��     �                                                                                      ����� ���?��     ��  8  '��{w� i  htw�����     ����� ���?��     �                         �������������������������������                              ����� ���?��     �����������@����������   	�0     ����� ���?��     �                                                                                      �   � ����      ����.z����>����� 0P  sv?�  ��     �   � ����      �                         �������������������������������                              �   � ����      �х\g!�DD0�ϯ���������0     �   � ����      �                                                     �@                              �   � ����      ��� V %�_{���� �`G��������     �   � ����      �                         �������������������������������                              �   � ����      ����������"#��?����D@   �p     �   � ����      �                                                                                      ����� ��?�      ���� ;��`��~    � �  ?�����     ����� ��?�      �                         �������������������������������                              ����� ��?�      ��<����q��"�����]�k����  ��     ����� ��?�      �                                                                                      ����� ��?�                                         ����� ��?�      �                                                                                    ����� ��?�      �������������������������������     ����� ��?�      �                                                                                      ����� �?����                                         ����� �?����     �                                                                                      ����� �?����                                         ����� �?����     �                                                                                      ����� ?�?����                                         ����� ?�?����     �                                                                                      ����� ?�?����                                         ����� ?�?����     �                                                                                      �   � ?�?���       �   x � �   x � �         �   � ?�?���     �                                                                                      �   � ?�?���       �   x � �   x � �         �   � ?�?���     �                                                                                      �   � ? ?���       �   x � �   x � �         �   � ? ?���     �                                                                                      �   � ? ?���       �   x � �   x � �         �   � ? ?���     �                                                                                      ����� ?             �   x � �   x � �         ����� ?           �                                                                                      ����� ?             �   x � �   x � �         ����� ?           �                                                                                      ����� >             �   x � �   x � �         ����� >           �                                                                                      ����� >             �   x � �   x � �         ����� >           �                                                                                      �����  �����        �   x � �   x � �         �����  �����      �                                                                                      �����  �����        �   x � �   x � �         �����  �����      �                                                                                      �����  �����        �   x � �   x � �         �����  �����      �                                                                                      �����  �����        �   x � �   x � �         �����  �����      �                                                                                       ��   �����        �   x � �   x � �          ��   �����      �                                                                                       ��   �����        �   x � �   x � �          ��   �����      �                                                                                       ��   �����        �   x � �   x � �          ��   �����      �                                                                                       ��   �����        �   x � �   x � �          ��   �����      �                                                                                       ��   � �        �   x � �   x � �          ��   � �      �                                                                                       ��   � �        �   x � �   x � �          ��   � �      �                                                                                       ��   � �        �   x � �   x � �          ��   � �      �                                                                                       ��   � �        �   x � �   x � �          ��   � �      �                                                                                    ������� � �        �   x � �   x � �       ������� � �      �                                                                                    ������� � �        �   x � �   x � �       ������� � �      �                                                                                    ������� � �        �   x � �   x � �       ������� � �      �                                                                                    ������� � �        �   x � �   x � �       ������� � �      �                                                                                    ������� � �        �   x � �   x � �       ������� � �      �                                                                                    ������� � �        �   x � �   x � �       ������� � �      �                                                                                    ������� � �        �   x � �   x � �       ������� � �      �                                                                                    ������� � �        �   x � �   x � �       ������� � �      �                                                                                      ��   � �        �   x � �   x � �         ��   � �      �                                                                                      ��   � �        �   x � �   x � �         ��   � �      �                                                                                      ��   � �        �   x � �   x � �         ��   � �      �                                                                                      ��   � �        �   x � �   x � �         ��   � �      �                                                                                      ��   � �        �   x � �   x � �         ��   � �      �                                                                                      ��   � �        �   x � �   x � �         ��   � �      �                                                                                      ��   � �        �   x � �   x � �         ��   � �      �                                                                                      ��   � �        �   x � �   x � �         ��   � �      �                                                                                                        �������������������������������                       �                                                                                                        �������������������������������                       �                                                                                                        �                                                    �                                                                                                        �                                                    �                                                                                                        �                                                    �                                                                                                        �                                                    �                                                                                                        �                                                    �                                                                                                        �                                                    �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            