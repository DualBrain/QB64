�P   ˀ�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 �������������������������������������������������������������������������������                                                                                �������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                              �������������������������������������������������������������������������������                                                                                �������������������������������������������������������������������������������                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                      � �   �                                             � �   �         �                                                                                      � �   �                                             � �   �         �                                                                                     � �   �                                            � �   �         �                                                                                     � �   �                                            � �   �         �                                                                                     � �   � ��                                         � �   � ��      �                                                                                     � �   � ��                                         � �   � ��      �                                     x       �� ��                                 � �   � ��                  0       ! �        � �   � ��      �                                                                                     � �   � ��                  x       �� �p        � �   � ��      �                             ?���   �    ������  ��                            �����������          ?���   �    ���� ��  ��   �����������      �                                                                                     �����������       >   ?���    �    ������  ��   �����������      �                          �   ����   �    ������  ��                            �����������          ����   �    ?���� ��  ��   �����������      �                                                                                     �����������       �   ���   �    ������  ��   �����������      �                         ��  �����  �   �������  ?��                            ����������<      �   �����  �    ����� ��  ��   ����������<      �                                                                                     ����������<      ��  �����  �   �������  ?��   ����������<      �                         ��  �����  �   �������  ��                            ����������<      ��  �����  �   ����� ��  ��   ����������<      �                                                                                     ����������<      ��  �����  �   �������  ��   ����������<      �                         ��  �����  �   �������  ���                            ?��?�� ���<     ��  ����  �   �������  ���   ?��?�� ���<     �                                                                                     ?��?�� ���<     ��  �����  ?�   ����� ��  ���   ?��?�� ���<     �                         ?��  ����  ���  ����� �� ���                            ?���� ���<?     ��  ���  ��  ����� ��  ��   ?���� ���<?     �                                                                                     ?���� ���<?     ?��  ����  ��   ����� �� ���   ?���� ���<?     �                         ?��  ����  ���  ����� �� ��                             ���� ����<|     ?��  ���  ���  ����� �� ��    ���� ����<|     �                                                                                     ���� ����<|     ?��  ����  ���  ?��|�� �� ��    ���� ����<|     �                         ?��  ����  ���  �� �� �� ��                             ����� ����<�     ��  ���  ��  �� �� �� ��    ����� ����<�     �                                                                                     ����� ����<�     ?��  ����  ���  �� �� �� ��    ����� ����<�     �                         ��  ����  ��  ��  �� �� ��                             � �   ����?�     ��  ���  ��  ��  �� �� ��    � �   ����?�     �                                                                                     � �   ����?�     ��  �� ��  ��  ��  �� �� ��    � �   ����?�     �                         ��  �� ��  �� ��  �� �� ��                             � �   ����?�     ��  � ��  ��  ��  �� �� ��    � �   ����?�     �                                                                                     � �   ����?�     ��  �� ��  ?�� ��  �� �� ��    � �   ����?�     �                         ��  �� ��  ?�� ��  �� �� ��                             ������ ����     ��  � ��  �� ��  �� �� ��    ������ ����     �                                                                                     ������ ����     ��  �� �  ?�� ��  �� �� ��    ������ ����     �                         ��  �� �  �� ��  �� �� ��                             ������ ����     ��  � �  �� ��  �� �� ��    ������ ����     �                                                                                     ������ ����     ��  �� �  �� ��  �� �� ��    ������ ����     �                         ��  �� �  �� ��  �� �� ��                              ����� ����        ��  �� �  �� ��  �� �� ��     ����� ����        �                                                                                      ����� ����        ��  � �  �� ��  �� �� ��     ����� ����        �                         ��  � ��  ?�� ��  �� �� ��                              ����� ����        ��  � ��  �� ��  �� �� ��     ����� ����        �                                                                                      ����� ����        ��  � �  ?�� ��  �� �� ��     ����� ����        �                         ��� � ��  ?�� ��  �� �� ��                              �   � �������     ��� � ��  ?�� ��  �� �� ��     �   � �������     �                                                                                      �   � �������     ��  � ��  ?�� ��  �� �� ��     �   � �������     �                         ��� ���  �� ��  �� �� ��                              �   � �������     ��� ���  �� ��  �� �� ��     �   � �������     �                                                                                      �   � �������     ��� � ��  �� ��  �� �� ��     �   � �������     �                         ?��� ���  ��� ��  �� �� ��                              �   � ������     ?��� ���  ��� ��  �� �� ��     �   � ������     �                         ?��� ���  ��� ��  �� �� ��                              �   � ������                                         �   � ������     �                         ?��� ���  ��� ��  �� �� ��                              �   � ������     ?��� ���  ��� ��  �� �� ��     �   � ������     �                                                                                      �   � ������     ?��� ���  ��� ��  �� �� ��     �   � ������     �                         ��� ��� ������  �� �� ��                              ����� ���<�     ��� ��� ������  �� �� ��     ����� ���<�     �                                                                                      ����� ���<�     ��� ��� ������  �� �� ��     ����� ���<�     �                         ���� ���� ������  �� �� ��                              ����� ���<�     ���� ���� ������  �� �� ��     ����� ���<�     �                                                                                      ����� ���<�     ��� ���  ������  �� �� ��     ����� ���<�     �                         ���� ���  �����  �� �� ��                              ����� ���?��     ���� ���  �����  �� �� ��     ����� ���?��     �                         ���� ���  �����  �� �� ��                              ����� ���?��     ���� ���  �����  �� �� ��     ����� ���?��     �                        ���� ���� �����  �� �� ��                              ����� ���?��     ���� ���� �����  �� �� ��     ����� ���?��     �                                                                                      ����� ���?��    ���� ���� �?����  �� �� ��     ����� ���?��     �                        ���� ���� �?����  �� �� ��                              �   � ����     ��� ���� �?����  �� �� ��     �   � ����      �                                                                                      �   � ����     ���� ���� �?����  �� �� ��     �   � ����      �                        ��� ���� �?����  �� �� ��                              �   � ����     ��� ���� �?����  �� �� ��     �   � ����      �                                                                                      �   � ����     ��� ���� �����  �� �� ��     �   � ����      �                        ��� ���� �����  �� �� ��                              ����� ��?�     ��� ���� �����  �� �� ��     ����� ��?�      �                        ��� ���� �����  �� �� ��                              ����� ��?�     ��� ���� �����  �� �� ��     ����� ��?�      �                        ��� ��� ?�����  �� �� ��                              ����� ��?�     ��� ��� ?�����  �� �� ��     ����� ��?�      �                                                                                      ����� ��?�     ��� ��� �����  �� �� ��     ����� ��?�      �                        �������� ?������  �� �� ��                              ����� �?����    �������� ?�����  �� �� ��     ����� �?����     �                                                                                      ����� �?����    ���� ��� ?������  �� �� ��     ����� �?����     �                        �������� ������  �� �� ��                              ����� ?�?����    �������� ?������  �� �� ��     ����� ?�?����     �                                                                                      ����� ?�?����    ������ �� ������  �� �� ��     ����� ?�?����     �                        ?������ �� �������  �� �� ��                              �   � ?�?���    ?������ �� �������  �� �� ��     �   � ?�?���     �                        ?������ �� �������  �� �� ��                              �   � ?�?���                                         �   � ?�?���     �                        ?������ � ��������  �� �� ��                              �   � ? ?���    ?����� � ��������  �� �� ��     �   � ? ?���     �                                                                                      �   � ? ?���    ?������ � �������  �� �� ��     �   � ? ?���     �                        ����� ���������  �� �� ��                              ����� ?          ?����� � ��������  �� �� ��     ����� ?           �                                                                                      ����� ?          ����� ?���������  �� �� ��     ����� ?           �                        ������� ?���������� �� �� ��                              ����� >          ���?���� ?��?������� �� �� ��     ����� >           �                                                                                      ����� >          ����� ?���������� �� �� ��     ����� >           �                        �������� ?���������� ���� ��                              �����  �����     ������� ?��������� ���� ��     �����  �����      �                                                                                      �����  �����     �������� ?���������� �� �� ��     �����  �����      �                       �������� ��������������� ��                              �����  �����     ������� ?��������������� ��     �����  �����      �                                                                                      �����  �����    �������� ������������� ��     �����  �����      �                       �������� ���������������� ��                               ��   �����    ������� ���������������� ��      ��   �����      �                                                                                       ��   �����    �������� ��������������� ��      ��   �����      �                       �������� ����������������� ?��                               ��   �����    ������� ����������������� ��      ��   �����      �                                                                                       ��   �����    �������� ���������������� ?��      ��   �����      �                       ������������������������� ��                               ��   � �    ����������������������� ��      ��   � �      �                                                                                       ��   � �    ������� ����������������� ?��      ��   � �      �                       �?��������?������������� ���                               ��   � �    �?�������?������������� ��       ��   � �      �                                                                                       ��   � �    �?��������������������� ��      ��   � �      �                       ��������?����?����������                             ������� � �    �������?�?���?����������    ������� � �      �                                                                                    ������� � �    ��������?����?��������s��    ������� � �      �                       ���������?�?�������������                             ������� � �    ���������?��������������    ������� � �      �                                                                                    ������� � �    ���������?�?�������������    ������� � �      �                       ���������?��������������                             ������� � �    ������������ ��� �������    ������� � �      �                                                                                    ������� � �    ���������?��������������    ������� � �      �                       ������������ ��� �������                             ������� � �    �� ���������� ��� �������    ������� � �      �                                                                                    ������� � �    ������������ ��� �����?��    ������� � �      �                       � � ����������  ��� ����?��                               ��   � �    � � ����������  �� ?����?��      ��   � �      �                                                                                      ��   � �    � � � ��� ���  ��� ����?��      ��   � �      �                       �   � ��� �  �  �� �����                               ��   � �    �   ~ ��� �  �  �� �����      ��   � �      �                                                                                      ��   � �    �   � ?��� �  �  �� � ���       ��   � �      �                       �   |      �  �                                             ��   � �    �   |         �                    ��   � �      �                                                                                      ��   � �    �   |      �  �                    ��   � �      �                       �   x         �                                             ��   � �    �   x         �                    ��   � �      �                                                                                      ��   � �    �   8          �                    ��   � �      �                                                                                                                                                              �                                                                                                                                                              �                                     B     @                                                                        B     @                                   �                                                                                                                    B     @                                   �                                     �                                                                              �                                         �                                                                                                                    �                                         �                                     �                                                                              �                                         �                                                                                                                    �                                         �                                     �s�,q�                                                                         �s�,q�                                    �                                                                                                                    �s�,q�                                    �                                     �
 ��Q                                                                         �
 ��Q                                    �                                                                                                                    �
 ��Q                                    �                                     �z'��                                                                         �z'��                                    �                                                                                                                    �z'��                                    �                                     ��(���                                                                         ��(���                                    �                                                                                                                    ��(���                                    �                                     ��(��Q                                                                         ��(��Q                                    �                                                                                                                    ��(��Q                                    �                                     �{Ǣq�                                                                         �{Ǣq�                                    �                                                                                                                    �{Ǣq�                                    �                                     �                                                                             �                                        �                                                                                                                    �                                        �                                     @    @                                                                        @    @                                   �                                                                                                                    @    @                                   �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                        �������������������������������                       �                                                                                                        �������������������������������                       �                                                                                                        �                                                    �                                                                                                        �                                                    �                                                                                                        �                                                    �                                                                                                        �                                                    �                                                                                                        �                                                    �                                                                                                        �                                                    �                                                                                                        �                                                    �                                                                                                        �                                                    �                          >|��                     ���                                                 �>|��                     ���                       �                          >|��                     ���                                                 �                                                    �                          !A                     P�                                                  �!A                     P�                        �                          !A                     P�                                                  �                                                    �                          !A                     P�                                                  �!A                     P�                        �                          !A                     P�                                                  �                                                    �                          !A                     P�                                                  �!A                     P�                        �                          !A                     P�                                                  �                                                    �                          >x�                     P�                                                  �>x�                     P�                        �                          >x�                     P�                                                  �                                                    �                          !@                     P�                                                  �!@                     P�                        �                          !@                     P�                                                  �                                                    �                          !@                     	P�                                                  �!@                     	P�                        �                          !@                     	P�                                                  �                                                    �                          !A                     Т                                                  �!A                     Т                        �                          !A                     Т                                                  �                                                    �                          !|��                     �"                                                  �!|��                     �"                        �                          !|��                     �"                                                  �                                                    �                                                    @                                                   �                          @                         �                                                    @                                                   �                                                    �                                                                                                        �                                                    �                                                                                                        �                                                    �                                                                                                        �                                                    �                                                                                                        �                                                    �                                                                                                        �                                                    �                                                                                                        �                                                    �                                                                                                        �������������������������������                       �                                                                                                        �������������������������������                       �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                                                                                                                                                              �                         ��                          ��                                                ��                          ��                       �                         �������������������������������                                                ��                          ��                       �                                                                                                        �������� |b��� �  �-�'f����                       �                         �������������������������������                                                ��    ����Y@ �� ����*ؙ?���                       �                                                                                                        �������   ���������s� �JA~p                       �                         �����������������������������~p                                                ��    ����EU@��!�������                       �                                                                                                        ��������|D��� ����  4Y���                       �                         ������������������������������                                                ��      SY@8��� A��˦^n|0                       �                                                                                                        ������    ݿ������   P����                       �                         �������������������������������                                                ��   ?�����"@@   _����Kg�2��0                       �                                                      @                                                �  �� vټ�C~�����  �,�'��                       �                         �������������������������������                                                ���� ���&C4���?� B��M�e���p                       �                                                                                                        ��������d� y��� }�wƱ``s�                       �                         �������������������������������                                                ��      �z���?����9N����                       �                                                                                      � �   �         ������ h�5�t#�  z w�9EEA�p     � �   �         �                         ������������������������������p                              � �   �         �� � ����~��������(ƺﺾ��     � �   �         �                          �                                                          � �   �         ��    �J�  c��   � 	� 1(}�    � �   �         �                         �������������������������������                             � �   �         ������� �:����?�����[����׾p    � �   �         �                                                                                     � �   � ��      �������  �]�?�� {��d9E��SA��    � �   � ��      �                         �������������������������������                             � �   � ��      ��   ����S�!�?���!�ƺi?��?p    � �   � ��      �                                                                                     � �   � ��      �8 ~  ?���]0 ���` ��D��    � �   � ��      �                         �?�����������������������������                             � �   � ��      ������� n��*�����p�/����k��0p    � �   � ��      �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            